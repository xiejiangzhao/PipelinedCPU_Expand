module InstRom
(
	input [3:0] addr,
	output [31:0] data
);
reg [31:0] ram [15:0];
always
	begin
		ram[0]=32'b000000_00011_00001_00010_00000_100000;//add  $2,$3,$1
		ram[1]=32'b000000_00011_00010_00010_00000_100010;//sub  $2,$3,$2
		ram[2]=32'b011100_00011_00000_00010_00000_100000;//clz   $2,$3
		ram[3]=32'b000000_00000_00001_00010_00000_000100;//sllv 
		ram[4]=32'b000000_00000_00001_00010_00100_000011;//sra
		ram[5]=32'b001010_00000_00010_0000_0000_1000_0000;//slti
		ram[6]=32'b001000_00000_00010_0000_0000_0000_1000;//addi
		ram[7]=32'b100011_00000_00010_0000_0000_0000_0100;//lw
		ram[8]=32'b010010_00000_00010_0000_0000_0000_0010;//lwl
		ram[9]=32'b010010_00000_00010_0000_0000_0000_0011;//lwl
		ram[10]=32'b010110_00000_00010_0000_0000_0000_0010;//lwr
		ram[11]=32'b101011_00000_00010_0000_0000_0011_0000;//sw
		ram[12]=32'b000110_00001_00000_0000_0000_0000_1000;//blez   $1
		ram[13]=32'b000010_00000_00000_0000_0000_0000_0010;//j        2
		ram[14]=32'b000000_00011_00001_00010_00000_100000;//add    $2,$3,$1
		//ram[15]=32'b000000_00011_00001_00010_00000_100000;//add    $2,$3,$1
	end
assign data = ram[addr];
endmodule
